`timescale 1ns / 100ps

module red_pitaya (
  input wire [1:1] adc_clk_i,
  output wire[7:0] led_o
);

  wire clk;
  assign clk = adc_clk_i[1];

  reg [128:0] counter;
  //assign led_o = counter[31:24];

  always @(posedge clk) begin
    counter <= counter + 1;
  end

  reg RST_N;
  initial begin
    RST_N = 0;
  end

  always @(posedge clk) begin
    RST_N <= counter > 1024 ? 1 : 0;
  end

  wire slave1_arready;
  wire slave1_rvalid;
  wire [11:0] slave1_rid;
  wire [31:0] slave1_rdata;
  wire [1:0] slave1_rresp;
  wire slave1_rlast;
  wire slave1_awready;
  wire slave1_wready;
  wire slave1_bvalid;
  wire [1:0] slave1_bresp;
  wire [11:0] slave1_bid;
  wire slave1_arvalid;
  wire [11:0] slave1_arid;
  wire [31:0] slave1_araddr;
  wire [7:0] slave1_arlen;
  wire [2:0] slave1_arsize;
  wire [1:0] slave1_arburst;
  wire slave1_arlock;
  wire [3:0] slave1_arcache;
  wire [2:0] slave1_arprot;
  wire [3:0] slave1_arqos;
  wire [3:0] slave1_arregion;
  wire slave1_rready;
  wire slave1_awvalid;
  wire [11:0] slave1_awid;
  wire [31:0] slave1_awaddr;
  wire [7:0] slave1_awlen;
  wire [2:0] slave1_awsize;
  wire [1:0] slave1_awburst;
  wire slave1_awlock;
  wire [3:0] slave1_awcache;
  wire [2:0] slave1_awprot;
  wire [3:0] slave1_awqos;
  wire [3:0] slave1_awregion;
  wire slave1_wvalid;
  wire [31:0] slave1_wdata;
  wire [3:0] slave1_wstrb;
  wire slave1_wlast;
  wire slave1_bready;

  wire slave0_arready;
  wire slave0_rvalid;
  wire [11:0] slave0_rid;
  wire [31:0] slave0_rdata;
  wire [1:0] slave0_rresp;
  wire slave0_rlast;
  wire slave0_awready;
  wire slave0_wready;
  wire slave0_bvalid;
  wire [1:0] slave0_bresp;
  wire [11:0] slave0_bid;
  wire slave0_arvalid;
  wire [11:0] slave0_arid;
  wire [31:0] slave0_araddr;
  wire [7:0] slave0_arlen;
  wire [2:0] slave0_arsize;
  wire [1:0] slave0_arburst;
  wire slave0_arlock;
  wire [3:0] slave0_arcache;
  wire [2:0] slave0_arprot;
  wire [3:0] slave0_arqos;
  wire [3:0] slave0_arregion;
  wire slave0_rready;
  wire slave0_awvalid;
  wire [11:0] slave0_awid;
  wire [31:0] slave0_awaddr;
  wire [7:0] slave0_awlen;
  wire [2:0] slave0_awsize;
  wire [1:0] slave0_awburst;
  wire slave0_awlock;
  wire [3:0] slave0_awcache;
  wire [2:0] slave0_awprot;
  wire [3:0] slave0_awqos;
  wire [3:0] slave0_awregion;
  wire slave0_wvalid;
  wire [31:0] slave0_wdata;
  wire [3:0] slave0_wstrb;
  wire slave0_wlast;
  wire slave0_bready;

  wire master0_arready;
  wire master0_rvalid;
  wire [2:0] master0_rid;
  wire [63:0] master0_rdata;
  wire [1:0] master0_rresp;
  wire master0_rlast;
  wire master0_awready;
  wire master0_wready;
  wire master0_bvalid;
  wire [1:0] master0_bresp;
  wire [2:0] master0_bid;
  wire master0_arvalid;
  wire [2:0] master0_arid;
  wire [31:0] master0_araddr;
  wire [7:0] master0_arlen;
  wire [2:0] master0_arsize;
  wire [1:0] master0_arburst;
  wire master0_arlock;
  wire [3:0] master0_arcache;
  wire [2:0] master0_arprot;
  wire [3:0] master0_arqos;
  wire [3:0] master0_arregion;
  wire master0_rready;
  wire master0_awvalid;
  wire [2:0] master0_awid;
  wire [31:0] master0_awaddr;
  wire [7:0] master0_awlen;
  wire [2:0] master0_awsize;
  wire [1:0] master0_awburst;
  wire master0_awlock;
  wire [3:0] master0_awcache;
  wire [2:0] master0_awprot;
  wire [3:0] master0_awqos;
  wire [3:0] master0_awregion;
  wire master0_wvalid;
  wire [63:0] master0_wdata;
  wire [7:0] master0_wstrb;
  wire master0_wlast;
  wire master0_bready;
  wire [4:0] master0_ruser;
  wire [4:0] master0_buser;
  wire [4:0] master0_wuser;
  wire [4:0] master0_aruser;
  wire [4:0] master0_awuser;

  mkSoc soc (
    .RST_N(RST_N),
    .CLK(clk),

    // Debug led
    .leds(led_o),

    // Slave interfaces
    .slave0_arready    (slave0_arready ),
    .slave0_rvalid     (slave0_rvalid  ),
    .slave0_rid        (slave0_rid     ),
    .slave0_rdata      (slave0_rdata   ),
    .slave0_rresp      (slave0_rresp   ),
    .slave0_rlast      (slave0_rlast   ),
    .slave0_awready    (slave0_awready ),
    .slave0_wready     (slave0_wready  ),
    .slave0_bvalid     (slave0_bvalid  ),
    .slave0_bresp      (slave0_bresp   ),
    .slave0_bid        (slave0_bid     ),
    .slave0_arvalid    (slave0_arvalid ),
    .slave0_arid       (slave0_arid    ),
    .slave0_araddr     (slave0_araddr  ),
    .slave0_arlen      (slave0_arlen   ),
    .slave0_arsize     (slave0_arsize  ),
    .slave0_arburst    (slave0_arburst ),
    .slave0_arlock     (slave0_arlock  ),
    .slave0_arcache    (slave0_arcache ),
    .slave0_arprot     (slave0_arprot  ),
    .slave0_arqos      (slave0_arqos   ),
    .slave0_arregion   (slave0_arregion),
    .slave0_rready     (slave0_rready  ),
    .slave0_awvalid    (slave0_awvalid ),
    .slave0_awid       (slave0_awid    ),
    .slave0_awaddr     (slave0_awaddr  ),
    .slave0_awlen      (slave0_awlen   ),
    .slave0_awsize     (slave0_awsize  ),
    .slave0_awburst    (slave0_awburst ),
    .slave0_awlock     (slave0_awlock  ),
    .slave0_awcache    (slave0_awcache ),
    .slave0_awprot     (slave0_awprot  ),
    .slave0_awqos      (slave0_awqos   ),
    .slave0_awregion   (slave0_awregion),
    .slave0_wvalid     (slave0_wvalid  ),
    .slave0_wdata      (slave0_wdata   ),
    .slave0_wstrb      (slave0_wstrb   ),
    .slave0_wlast      (slave0_wlast   ),
    .slave0_bready     (slave0_bready  ),

    .slave1_arready    (slave1_arready ),
    .slave1_rvalid     (slave1_rvalid  ),
    .slave1_rid        (slave1_rid     ),
    .slave1_rdata      (slave1_rdata   ),
    .slave1_rresp      (slave1_rresp   ),
    .slave1_rlast      (slave1_rlast   ),
    .slave1_awready    (slave1_awready ),
    .slave1_wready     (slave1_wready  ),
    .slave1_bvalid     (slave1_bvalid  ),
    .slave1_bresp      (slave1_bresp   ),
    .slave1_bid        (slave1_bid     ),
    .slave1_arvalid    (slave1_arvalid ),
    .slave1_arid       (slave1_arid    ),
    .slave1_araddr     (slave1_araddr  ),
    .slave1_arlen      (slave1_arlen   ),
    .slave1_arsize     (slave1_arsize  ),
    .slave1_arburst    (slave1_arburst ),
    .slave1_arlock     (slave1_arlock  ),
    .slave1_arcache    (slave1_arcache ),
    .slave1_arprot     (slave1_arprot  ),
    .slave1_arqos      (slave1_arqos   ),
    .slave1_arregion   (slave1_arregion),
    .slave1_rready     (slave1_rready  ),
    .slave1_awvalid    (slave1_awvalid ),
    .slave1_awid       (slave1_awid    ),
    .slave1_awaddr     (slave1_awaddr  ),
    .slave1_awlen      (slave1_awlen   ),
    .slave1_awsize     (slave1_awsize  ),
    .slave1_awburst    (slave1_awburst ),
    .slave1_awlock     (slave1_awlock  ),
    .slave1_awcache    (slave1_awcache ),
    .slave1_awprot     (slave1_awprot  ),
    .slave1_awqos      (slave1_awqos   ),
    .slave1_awregion   (slave1_awregion),
    .slave1_wvalid     (slave1_wvalid  ),
    .slave1_wdata      (slave1_wdata   ),
    .slave1_wstrb      (slave1_wstrb   ),
    .slave1_wlast      (slave1_wlast   ),
    .slave1_bready     (slave1_bready  ),

    // Master interface
    .master0_arready    (master0_arready ),
    .master0_rvalid     (master0_rvalid  ),
    .master0_rid        (master0_rid     ),
    .master0_rdata      (master0_rdata   ),
    .master0_rresp      (master0_rresp   ),
    .master0_rlast      (master0_rlast   ),
    .master0_awready    (master0_awready ),
    .master0_wready     (master0_wready  ),
    .master0_bvalid     (master0_bvalid  ),
    .master0_bresp      (master0_bresp   ),
    .master0_bid        (master0_bid     ),
    .master0_arvalid    (master0_arvalid ),
    .master0_arid       (master0_arid    ),
    .master0_araddr     (master0_araddr  ),
    .master0_arlen      (master0_arlen   ),
    .master0_arsize     (master0_arsize  ),
    .master0_arburst    (master0_arburst ),
    .master0_arlock     (master0_arlock  ),
    .master0_arcache    (master0_arcache ),
    .master0_arprot     (master0_arprot  ),
    .master0_arqos      (master0_arqos   ),
    .master0_arregion   (master0_arregion),
    .master0_rready     (master0_rready  ),
    .master0_awvalid    (master0_awvalid ),
    .master0_awid       (master0_awid    ),
    .master0_awaddr     (master0_awaddr  ),
    .master0_awlen      (master0_awlen   ),
    .master0_awsize     (master0_awsize  ),
    .master0_awburst    (master0_awburst ),
    .master0_awlock     (master0_awlock  ),
    .master0_awcache    (master0_awcache ),
    .master0_awprot     (master0_awprot  ),
    .master0_awqos      (master0_awqos   ),
    .master0_awregion   (master0_awregion),
    .master0_wvalid     (master0_wvalid  ),
    .master0_wdata      (master0_wdata   ),
    .master0_wstrb      (master0_wstrb   ),
    .master0_wlast      (master0_wlast   ),
    .master0_bready     (master0_bready  ),
    .master0_ruser      (master0_ruser   ),
    .master0_buser      (master0_buser   ),
    .master0_aruser     (master0_aruser  ),
    .master0_wuser      (master0_wuser   ),
    .master0_awuser     (master0_awuser  )
  );

  //PS7 zynq7 ();

   PS7 zynq7 (
     .DMA0DATYPE(),
     .DMA0DAVALID(),
     .DMA0DRREADY(),
     .DMA0RSTN(),
     .DMA1DATYPE(),
     .DMA1DAVALID(),
     .DMA1DRREADY(),
     .DMA1RSTN(),
     .DMA2DATYPE(),
     .DMA2DAVALID(),
     .DMA2DRREADY(),
     .DMA2RSTN(),
     .DMA3DATYPE(),
     .DMA3DAVALID(),
     .DMA3DRREADY(),
     .DMA3RSTN(),
     .EMIOCAN0PHYTX(),
     .EMIOCAN1PHYTX(),
     .EMIOENET0GMIITXD(),
     .EMIOENET0GMIITXEN(),
     .EMIOENET0GMIITXER(),
     .EMIOENET0MDIOMDC(),
     .EMIOENET0MDIOO(),
     .EMIOENET0MDIOTN(),
     .EMIOENET0PTPDELAYREQRX(),
     .EMIOENET0PTPDELAYREQTX(),
     .EMIOENET0PTPPDELAYREQRX(),
     .EMIOENET0PTPPDELAYREQTX(),
     .EMIOENET0PTPPDELAYRESPRX(),
     .EMIOENET0PTPPDELAYRESPTX(),
     .EMIOENET0PTPSYNCFRAMERX(),
     .EMIOENET0PTPSYNCFRAMETX(),
     .EMIOENET0SOFRX(),
     .EMIOENET0SOFTX(),
     .EMIOENET1GMIITXD(),
     .EMIOENET1GMIITXEN(),
     .EMIOENET1GMIITXER(),
     .EMIOENET1MDIOMDC(),
     .EMIOENET1MDIOO(),
     .EMIOENET1MDIOTN(),
     .EMIOENET1PTPDELAYREQRX(),
     .EMIOENET1PTPDELAYREQTX(),
     .EMIOENET1PTPPDELAYREQRX(),
     .EMIOENET1PTPPDELAYREQTX(),
     .EMIOENET1PTPPDELAYRESPRX(),
     .EMIOENET1PTPPDELAYRESPTX(),
     .EMIOENET1PTPSYNCFRAMERX(),
     .EMIOENET1PTPSYNCFRAMETX(),
     .EMIOENET1SOFRX(),
     .EMIOENET1SOFTX(),
     .EMIOGPIOO(),
     .EMIOGPIOTN(),
     .EMIOI2C0SCLO(),
     .EMIOI2C0SCLTN(),
     .EMIOI2C0SDAO(),
     .EMIOI2C0SDATN(),
     .EMIOI2C1SCLO(),
     .EMIOI2C1SCLTN(),
     .EMIOI2C1SDAO(),
     .EMIOI2C1SDATN(),
     .EMIOPJTAGTDO(),
     .EMIOPJTAGTDTN(),
     .EMIOSDIO0BUSPOW(),
     .EMIOSDIO0BUSVOLT(),
     .EMIOSDIO0CLK(),
     .EMIOSDIO0CMDO(),
     .EMIOSDIO0CMDTN(),
     .EMIOSDIO0DATAO(),
     .EMIOSDIO0DATATN(),
     .EMIOSDIO0LED(),
     .EMIOSDIO1BUSPOW(),
     .EMIOSDIO1BUSVOLT(),
     .EMIOSDIO1CLK(),
     .EMIOSDIO1CMDO(),
     .EMIOSDIO1CMDTN(),
     .EMIOSDIO1DATAO(),
     .EMIOSDIO1DATATN(),
     .EMIOSDIO1LED(),
     .EMIOSPI0MO(),
     .EMIOSPI0MOTN(),
     .EMIOSPI0SCLKO(),
     .EMIOSPI0SCLKTN(),
     .EMIOSPI0SO(),
     .EMIOSPI0SSNTN(),
     .EMIOSPI0SSON(),
     .EMIOSPI0STN(),
     .EMIOSPI1MO(),
     .EMIOSPI1MOTN(),
     .EMIOSPI1SCLKO(),
     .EMIOSPI1SCLKTN(),
     .EMIOSPI1SO(),
     .EMIOSPI1SSNTN(),
     .EMIOSPI1SSON(),
     .EMIOSPI1STN(),
     .EMIOTRACECTL(),
     .EMIOTRACEDATA(),
     .EMIOTTC0WAVEO(),
     .EMIOTTC1WAVEO(),
     .EMIOUART0DTRN(),
     .EMIOUART0RTSN(),
     .EMIOUART0TX(),
     .EMIOUART1DTRN(),
     .EMIOUART1RTSN(),
     .EMIOUART1TX(),
     .EMIOUSB0PORTINDCTL(),
     .EMIOUSB0VBUSPWRSELECT(),
     .EMIOUSB1PORTINDCTL(),
     .EMIOUSB1VBUSPWRSELECT(),
     .EMIOWDTRSTO(),
     .EVENTEVENTO(),
     .EVENTSTANDBYWFE(),
     .EVENTSTANDBYWFI(),
     .FCLKCLK(),
     .FCLKRESETN(),
     .FTMTF2PTRIGACK(),
     .FTMTP2FDEBUG(),
     .FTMTP2FTRIG(),
     .IRQP2F(),
     .MAXIGP0ARADDR(slave0_araddr),
     .MAXIGP0ARBURST(slave0_arburst),
     .MAXIGP0ARCACHE(slave0_arcache),
     .MAXIGP0ARESETN(),
     .MAXIGP0ARID(slave0_arid),
     .MAXIGP0ARLEN(slave0_arlen),
     .MAXIGP0ARLOCK(slave0_arlock),
     .MAXIGP0ARPROT(slave0_arprot),
     .MAXIGP0ARQOS(slave0_arqos),
     .MAXIGP0ARSIZE(slave0_arsize),
     .MAXIGP0ARVALID(slave0_arvalid),
     .MAXIGP0AWADDR(slave0_awaddr),
     .MAXIGP0AWBURST(slave0_awburst),
     .MAXIGP0AWCACHE(slave0_awcache),
     .MAXIGP0AWID(slave0_awid),
     .MAXIGP0AWLEN(slave0_awlen),
     .MAXIGP0AWLOCK(slave0_awlock),
     .MAXIGP0AWPROT(slave0_awprot),
     .MAXIGP0AWQOS(slave0_awqos),
     .MAXIGP0AWSIZE(slave0_awsize),
     .MAXIGP0AWVALID(slave0_awvalid),
     .MAXIGP0BREADY(slave0_bready),
     .MAXIGP0RREADY(slave0_rready),
     .MAXIGP0WDATA(slave0_wdata),
     .MAXIGP0WID(),
     .MAXIGP0WLAST(slave0_wlast),
     .MAXIGP0WSTRB(slave0_wstrb),
     .MAXIGP0WVALID(slave0_wvalid),
     .MAXIGP1ARADDR(slave1_araddr),
     .MAXIGP1ARBURST(slave1_arburst),
     .MAXIGP1ARCACHE(slave1_arcache),
     .MAXIGP1ARESETN(),
     .MAXIGP1ARID(slave1_arid),
     .MAXIGP1ARLEN(slave1_arlen),
     .MAXIGP1ARLOCK(slave1_arlock),
     .MAXIGP1ARPROT(slave1_arprot),
     .MAXIGP1ARQOS(slave1_arqos),
     .MAXIGP1ARSIZE(slave1_arsize),
     .MAXIGP1ARVALID(slave1_arvalid),
     .MAXIGP1AWADDR(slave1_awaddr),
     .MAXIGP1AWBURST(slave1_awburst),
     .MAXIGP1AWCACHE(slave1_awcache),
     .MAXIGP1AWID(slave1_awid),
     .MAXIGP1AWLEN(slave1_awlen),
     .MAXIGP1AWLOCK(slave1_awlock),
     .MAXIGP1AWPROT(slave1_awprot),
     .MAXIGP1AWQOS(slave1_awqos),
     .MAXIGP1AWSIZE(slave1_awsize),
     .MAXIGP1AWVALID(slave1_awvalid),
     .MAXIGP1BREADY(slave1_bready),
     .MAXIGP1RREADY(slave1_rready),
     .MAXIGP1WDATA(slave1_wdata),
     .MAXIGP1WID(),
     .MAXIGP1WLAST(slave1_wlast),
     .MAXIGP1WSTRB(slave1_wstrb),
     .MAXIGP1WVALID(slave1_wvalid),
     .SAXIACPARESETN(),
     .SAXIACPARREADY(),
     .SAXIACPAWREADY(),
     .SAXIACPBID(),
     .SAXIACPBRESP(),
     .SAXIACPBVALID(),
     .SAXIACPRDATA(),
     .SAXIACPRID(),
     .SAXIACPRLAST(),
     .SAXIACPRRESP(),
     .SAXIACPRVALID(),
     .SAXIACPWREADY(),
     .SAXIGP0ARESETN(),
     .SAXIGP0ARREADY(),
     .SAXIGP0AWREADY(),
     .SAXIGP0BID(),
     .SAXIGP0BRESP(),
     .SAXIGP0BVALID(),
     .SAXIGP0RDATA(),
     .SAXIGP0RID(),
     .SAXIGP0RLAST(),
     .SAXIGP0RRESP(),
     .SAXIGP0RVALID(),
     .SAXIGP0WREADY(),
     .SAXIGP1ARESETN(),
     .SAXIGP1ARREADY(),
     .SAXIGP1AWREADY(),
     .SAXIGP1BID(),
     .SAXIGP1BRESP(),
     .SAXIGP1BVALID(),
     .SAXIGP1RDATA(),
     .SAXIGP1RID(),
     .SAXIGP1RLAST(),
     .SAXIGP1RRESP(),
     .SAXIGP1RVALID(),
     .SAXIGP1WREADY(),
     .SAXIHP0ARESETN(),
     .SAXIHP0ARREADY(),
     .SAXIHP0AWREADY(),
     .SAXIHP0BID(),
     .SAXIHP0BRESP(),
     .SAXIHP0BVALID(),
     .SAXIHP0RACOUNT(),
     .SAXIHP0RCOUNT(),
     .SAXIHP0RDATA(),
     .SAXIHP0RID(),
     .SAXIHP0RLAST(),
     .SAXIHP0RRESP(),
     .SAXIHP0RVALID(),
     .SAXIHP0WACOUNT(),
     .SAXIHP0WCOUNT(),
     .SAXIHP0WREADY(),
     .SAXIHP1ARESETN(),
     .SAXIHP1ARREADY(),
     .SAXIHP1AWREADY(),
     .SAXIHP1BID(),
     .SAXIHP1BRESP(),
     .SAXIHP1BVALID(),
     .SAXIHP1RACOUNT(),
     .SAXIHP1RCOUNT(),
     .SAXIHP1RDATA(),
     .SAXIHP1RID(),
     .SAXIHP1RLAST(),
     .SAXIHP1RRESP(),
     .SAXIHP1RVALID(),
     .SAXIHP1WACOUNT(),
     .SAXIHP1WCOUNT(),
     .SAXIHP1WREADY(),
     .SAXIHP2ARESETN(),
     .SAXIHP2ARREADY(),
     .SAXIHP2AWREADY(),
     .SAXIHP2BID(),
     .SAXIHP2BRESP(),
     .SAXIHP2BVALID(),
     .SAXIHP2RACOUNT(),
     .SAXIHP2RCOUNT(),
     .SAXIHP2RDATA(),
     .SAXIHP2RID(),
     .SAXIHP2RLAST(),
     .SAXIHP2RRESP(),
     .SAXIHP2RVALID(),
     .SAXIHP2WACOUNT(),
     .SAXIHP2WCOUNT(),
     .SAXIHP2WREADY(),
     .SAXIHP3ARESETN(),
     .SAXIHP3ARREADY(),
     .SAXIHP3AWREADY(),
     .SAXIHP3BID(),
     .SAXIHP3BRESP(),
     .SAXIHP3BVALID(),
     .SAXIHP3RACOUNT(),
     .SAXIHP3RCOUNT(),
     .SAXIHP3RDATA(),
     .SAXIHP3RID(),
     .SAXIHP3RLAST(),
     .SAXIHP3RRESP(),
     .SAXIHP3RVALID(),
     .SAXIHP3WACOUNT(),
     .SAXIHP3WCOUNT(),
     .SAXIHP3WREADY(),
     .DDRA(),
     .DDRBA(),
     .DDRCASB(),
     .DDRCKE(),
     .DDRCKN(),
     .DDRCKP(),
     .DDRCSB(),
     .DDRDM(),
     .DDRDQ(),
     .DDRDQSN(),
     .DDRDQSP(),
     .DDRDRSTB(),
     .DDRODT(),
     .DDRRASB(),
     .DDRVRN(),
     .DDRVRP(),
     .DDRWEB(),
     .MIO(),
     .PSCLK(),
     .PSPORB(),
     .PSSRSTB(),
     .DDRARB(),
     .DMA0ACLK(),
     .DMA0DAREADY(),
     .DMA0DRLAST(),
     .DMA0DRTYPE(),
     .DMA0DRVALID(),
     .DMA1ACLK(),
     .DMA1DAREADY(),
     .DMA1DRLAST(),
     .DMA1DRTYPE(),
     .DMA1DRVALID(),
     .DMA2ACLK(),
     .DMA2DAREADY(),
     .DMA2DRLAST(),
     .DMA2DRTYPE(),
     .DMA2DRVALID(),
     .DMA3ACLK(),
     .DMA3DAREADY(),
     .DMA3DRLAST(),
     .DMA3DRTYPE(),
     .DMA3DRVALID(),
     .EMIOCAN0PHYRX(),
     .EMIOCAN1PHYRX(),
     .EMIOENET0EXTINTIN(),
     .EMIOENET0GMIICOL(),
     .EMIOENET0GMIICRS(),
     .EMIOENET0GMIIRXCLK(),
     .EMIOENET0GMIIRXD(),
     .EMIOENET0GMIIRXDV(),
     .EMIOENET0GMIIRXER(),
     .EMIOENET0GMIITXCLK(),
     .EMIOENET0MDIOI(),
     .EMIOENET1EXTINTIN(),
     .EMIOENET1GMIICOL(),
     .EMIOENET1GMIICRS(),
     .EMIOENET1GMIIRXCLK(),
     .EMIOENET1GMIIRXD(),
     .EMIOENET1GMIIRXDV(),
     .EMIOENET1GMIIRXER(),
     .EMIOENET1GMIITXCLK(),
     .EMIOENET1MDIOI(),
     .EMIOGPIOI(),
     .EMIOI2C0SCLI(),
     .EMIOI2C0SDAI(),
     .EMIOI2C1SCLI(),
     .EMIOI2C1SDAI(),
     .EMIOPJTAGTCK(),
     .EMIOPJTAGTDI(),
     .EMIOPJTAGTMS(),
     .EMIOSDIO0CDN(),
     .EMIOSDIO0CLKFB(),
     .EMIOSDIO0CMDI(),
     .EMIOSDIO0DATAI(),
     .EMIOSDIO0WP(),
     .EMIOSDIO1CDN(),
     .EMIOSDIO1CLKFB(),
     .EMIOSDIO1CMDI(),
     .EMIOSDIO1DATAI(),
     .EMIOSDIO1WP(),
     .EMIOSPI0MI(),
     .EMIOSPI0SCLKI(),
     .EMIOSPI0SI(),
     .EMIOSPI0SSIN(),
     .EMIOSPI1MI(),
     .EMIOSPI1SCLKI(),
     .EMIOSPI1SI(),
     .EMIOSPI1SSIN(),
     .EMIOSRAMINTIN(),
     .EMIOTRACECLK(),
     .EMIOTTC0CLKI(),
     .EMIOTTC1CLKI(),
     .EMIOUART0CTSN(),
     .EMIOUART0DCDN(),
     .EMIOUART0DSRN(),
     .EMIOUART0RIN(),
     .EMIOUART0RX(),
     .EMIOUART1CTSN(),
     .EMIOUART1DCDN(),
     .EMIOUART1DSRN(),
     .EMIOUART1RIN(),
     .EMIOUART1RX(),
     .EMIOUSB0VBUSPWRFAULT(),
     .EMIOUSB1VBUSPWRFAULT(),
     .EMIOWDTCLKI(),
     .EVENTEVENTI(),
     .FCLKCLKTRIGN(),
     .FPGAIDLEN(),
     .FTMDTRACEINATID(),
     .FTMDTRACEINCLOCK(),
     .FTMDTRACEINDATA(),
     .FTMDTRACEINVALID(),
     .FTMTF2PDEBUG(),
     .FTMTF2PTRIG(),
     .FTMTP2FTRIGACK(),
     .IRQF2P(),
     .MAXIGP0ACLK(clk),
     .MAXIGP0ARREADY(slave0_arready),
     .MAXIGP0AWREADY(slave0_awready),
     .MAXIGP0BID(slave0_bid),
     .MAXIGP0BRESP(slave0_bresp),
     .MAXIGP0BVALID(slave0_bvalid),
     .MAXIGP0RDATA(slave0_rdata),
     .MAXIGP0RID(slave0_rid),
     .MAXIGP0RLAST(slave0_rlast),
     .MAXIGP0RRESP(slave0_rresp),
     .MAXIGP0RVALID(slave0_rvalid),
     .MAXIGP0WREADY(slave0_wready),
     .MAXIGP1ACLK(clk),
     .MAXIGP1ARREADY(slave1_arready),
     .MAXIGP1AWREADY(slave1_awready),
     .MAXIGP1BID(slave1_bid),
     .MAXIGP1BRESP(slave1_bresp),
     .MAXIGP1BVALID(slave1_bvalid),
     .MAXIGP1RDATA(slave1_rdata),
     .MAXIGP1RID(slave1_rid),
     .MAXIGP1RLAST(slave1_rlast),
     .MAXIGP1RRESP(slave1_rresp),
     .MAXIGP1RVALID(slave1_rvalid),
     .MAXIGP1WREADY(slave1_wready),
     .SAXIACPACLK(),
     .SAXIACPARADDR(),
     .SAXIACPARBURST(),
     .SAXIACPARCACHE(),
     .SAXIACPARID(),
     .SAXIACPARLEN(),
     .SAXIACPARLOCK(),
     .SAXIACPARPROT(),
     .SAXIACPARQOS(),
     .SAXIACPARSIZE(),
     .SAXIACPARUSER(),
     .SAXIACPARVALID(),
     .SAXIACPAWADDR(),
     .SAXIACPAWBURST(),
     .SAXIACPAWCACHE(),
     .SAXIACPAWID(),
     .SAXIACPAWLEN(),
     .SAXIACPAWLOCK(),
     .SAXIACPAWPROT(),
     .SAXIACPAWQOS(),
     .SAXIACPAWSIZE(),
     .SAXIACPAWUSER(),
     .SAXIACPAWVALID(),
     .SAXIACPBREADY(),
     .SAXIACPRREADY(),
     .SAXIACPWDATA(),
     .SAXIACPWID(),
     .SAXIACPWLAST(),
     .SAXIACPWSTRB(),
     .SAXIACPWVALID(),
     .SAXIGP0ACLK(),
     .SAXIGP0ARADDR(),
     .SAXIGP0ARBURST(),
     .SAXIGP0ARCACHE(),
     .SAXIGP0ARID(),
     .SAXIGP0ARLEN(),
     .SAXIGP0ARLOCK(),
     .SAXIGP0ARPROT(),
     .SAXIGP0ARQOS(),
     .SAXIGP0ARSIZE(),
     .SAXIGP0ARVALID(),
     .SAXIGP0AWADDR(),
     .SAXIGP0AWBURST(),
     .SAXIGP0AWCACHE(),
     .SAXIGP0AWID(),
     .SAXIGP0AWLEN(),
     .SAXIGP0AWLOCK(),
     .SAXIGP0AWPROT(),
     .SAXIGP0AWQOS(),
     .SAXIGP0AWSIZE(),
     .SAXIGP0AWVALID(),
     .SAXIGP0BREADY(),
     .SAXIGP0RREADY(),
     .SAXIGP0WDATA(),
     .SAXIGP0WID(),
     .SAXIGP0WLAST(),
     .SAXIGP0WSTRB(),
     .SAXIGP0WVALID(),
     .SAXIGP1ACLK(),
     .SAXIGP1ARADDR(),
     .SAXIGP1ARBURST(),
     .SAXIGP1ARCACHE(),
     .SAXIGP1ARID(),
     .SAXIGP1ARLEN(),
     .SAXIGP1ARLOCK(),
     .SAXIGP1ARPROT(),
     .SAXIGP1ARQOS(),
     .SAXIGP1ARSIZE(),
     .SAXIGP1ARVALID(),
     .SAXIGP1AWADDR(),
     .SAXIGP1AWBURST(),
     .SAXIGP1AWCACHE(),
     .SAXIGP1AWID(),
     .SAXIGP1AWLEN(),
     .SAXIGP1AWLOCK(),
     .SAXIGP1AWPROT(),
     .SAXIGP1AWQOS(),
     .SAXIGP1AWSIZE(),
     .SAXIGP1AWVALID(),
     .SAXIGP1BREADY(),
     .SAXIGP1RREADY(),
     .SAXIGP1WDATA(),
     .SAXIGP1WID(),
     .SAXIGP1WLAST(),
     .SAXIGP1WSTRB(),
     .SAXIGP1WVALID(),
     .SAXIHP0ACLK(),
     .SAXIHP0ARADDR(),
     .SAXIHP0ARBURST(),
     .SAXIHP0ARCACHE(),
     .SAXIHP0ARID(),
     .SAXIHP0ARLEN(),
     .SAXIHP0ARLOCK(),
     .SAXIHP0ARPROT(),
     .SAXIHP0ARQOS(),
     .SAXIHP0ARSIZE(),
     .SAXIHP0ARVALID(),
     .SAXIHP0AWADDR(),
     .SAXIHP0AWBURST(),
     .SAXIHP0AWCACHE(),
     .SAXIHP0AWID(),
     .SAXIHP0AWLEN(),
     .SAXIHP0AWLOCK(),
     .SAXIHP0AWPROT(),
     .SAXIHP0AWQOS(),
     .SAXIHP0AWSIZE(),
     .SAXIHP0AWVALID(),
     .SAXIHP0BREADY(),
     .SAXIHP0RDISSUECAP1EN(),
     .SAXIHP0RREADY(),
     .SAXIHP0WDATA(),
     .SAXIHP0WID(),
     .SAXIHP0WLAST(),
     .SAXIHP0WRISSUECAP1EN(),
     .SAXIHP0WSTRB(),
     .SAXIHP0WVALID(),
     .SAXIHP1ACLK(),
     .SAXIHP1ARADDR(),
     .SAXIHP1ARBURST(),
     .SAXIHP1ARCACHE(),
     .SAXIHP1ARID(),
     .SAXIHP1ARLEN(),
     .SAXIHP1ARLOCK(),
     .SAXIHP1ARPROT(),
     .SAXIHP1ARQOS(),
     .SAXIHP1ARSIZE(),
     .SAXIHP1ARVALID(),
     .SAXIHP1AWADDR(),
     .SAXIHP1AWBURST(),
     .SAXIHP1AWCACHE(),
     .SAXIHP1AWID(),
     .SAXIHP1AWLEN(),
     .SAXIHP1AWLOCK(),
     .SAXIHP1AWPROT(),
     .SAXIHP1AWQOS(),
     .SAXIHP1AWSIZE(),
     .SAXIHP1AWVALID(),
     .SAXIHP1BREADY(),
     .SAXIHP1RDISSUECAP1EN(),
     .SAXIHP1RREADY(),
     .SAXIHP1WDATA(),
     .SAXIHP1WID(),
     .SAXIHP1WLAST(),
     .SAXIHP1WRISSUECAP1EN(),
     .SAXIHP1WSTRB(),
     .SAXIHP1WVALID(),
     .SAXIHP2ACLK(),
     .SAXIHP2ARADDR(),
     .SAXIHP2ARBURST(),
     .SAXIHP2ARCACHE(),
     .SAXIHP2ARID(),
     .SAXIHP2ARLEN(),
     .SAXIHP2ARLOCK(),
     .SAXIHP2ARPROT(),
     .SAXIHP2ARQOS(),
     .SAXIHP2ARSIZE(),
     .SAXIHP2ARVALID(),
     .SAXIHP2AWADDR(),
     .SAXIHP2AWBURST(),
     .SAXIHP2AWCACHE(),
     .SAXIHP2AWID(),
     .SAXIHP2AWLEN(),
     .SAXIHP2AWLOCK(),
     .SAXIHP2AWPROT(),
     .SAXIHP2AWQOS(),
     .SAXIHP2AWSIZE(),
     .SAXIHP2AWVALID(),
     .SAXIHP2BREADY(),
     .SAXIHP2RDISSUECAP1EN(),
     .SAXIHP2RREADY(),
     .SAXIHP2WDATA(),
     .SAXIHP2WID(),
     .SAXIHP2WLAST(),
     .SAXIHP2WRISSUECAP1EN(),
     .SAXIHP2WSTRB(),
     .SAXIHP2WVALID(),
     .SAXIHP3ACLK(),
     .SAXIHP3ARADDR(),
     .SAXIHP3ARBURST(),
     .SAXIHP3ARCACHE(),
     .SAXIHP3ARID(),
     .SAXIHP3ARLEN(),
     .SAXIHP3ARLOCK(),
     .SAXIHP3ARPROT(),
     .SAXIHP3ARQOS(),
     .SAXIHP3ARSIZE(),
     .SAXIHP3ARVALID(),
     .SAXIHP3AWADDR(),
     .SAXIHP3AWBURST(),
     .SAXIHP3AWCACHE(),
     .SAXIHP3AWID(),
     .SAXIHP3AWLEN(),
     .SAXIHP3AWLOCK(),
     .SAXIHP3AWPROT(),
     .SAXIHP3AWQOS(),
     .SAXIHP3AWSIZE(),
     .SAXIHP3AWVALID(),
     .SAXIHP3BREADY(),
     .SAXIHP3RDISSUECAP1EN(),
     .SAXIHP3RREADY(),
     .SAXIHP3WDATA(),
     .SAXIHP3WID(),
     .SAXIHP3WLAST(),
     .SAXIHP3WRISSUECAP1EN(),
     .SAXIHP3WSTRB(),
     .SAXIHP3WVALID()
 );
endmodule

